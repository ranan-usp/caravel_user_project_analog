** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/analog_switch.sch
**.subckt analog_switch IN control OUT
*.ipin IN
*.ipin control
*.opin OUT
x1 control OUT IN net1 transmission_gate
x2 control net1 not
**.ends

* expanding   symbol:  transmission_gate.sym # of pins=4
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/transmission_gate.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/transmission_gate.sch
.subckt transmission_gate  GP OUT IN GN
*.opin OUT
*.ipin IN
*.ipin GN
*.ipin GP
XM1 OUT GN IN GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT GP IN VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=3 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  not.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/not.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/not.sch
.subckt not  a y
*.ipin a
*.opin y
XM1 y a GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
