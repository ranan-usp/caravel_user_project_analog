** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/untitled.sch
**.subckt untitled
x1 vout en vdd vdd vss bootstrapped_sw_hv
V1 vdd GND 1.4
V2 vss GND 0
V3 en GND PULSE(0 1 10e-6 1e-9 1e-9 2e-6 4e-6)
C1 vout GND 1p m=1
V4 vdd GND vin
**** begin user architecture code

*.options method trap
*.options gmin 1e-15
*.options abstol 1e-15
*.options reltol 0.0001
*.options vntol 0.1e-6
*
*.include \$::DESIGN_PATH\/switches/bootstrapped_sw.sp

.param vin=0.7
.param MC_SWITCH=0

*.tran 100e-9 4e-6
.temp 85

.control
save all
tran 100e-9 16e-6 uic
run


* settle values
meas tran vset find v(vout) at=3.99e-6
meas tran vg_end find v(xsw.vg) at=3.99e-6
meas tran vin_end find v(vin) at=3.99e-6

let vgs_end=vg_end-vin_end

* max values
meas tran vg_max max xsw.vg
meas tran vs_max max xsw.vs
meas tran vbsl_max max xsw.vbsl
meas tran vbsh_max max xsw.vbsh

* min values
meas tran vg_min min xsw.vg
meas tran vs_min min xsw.vs
meas tran vbsl_min min xsw.vbsl
meas tran vbsh_min min xsw.vbsh


* print results
print vset
print vgs_end

print vg_max
print vs_max
print vbsl_max
print vbsh_max
print vg_min
print vs_min
print vbsl_min
print vbsh_min

.endc


 .lib /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice

**** end user architecture code
**.ends

* expanding   symbol:  adc/bootstrapped_sw_hv.sym # of pins=5
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/bootstrapped_sw_hv.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/bootstrapped_sw_hv.sch
.subckt bootstrapped_sw_hv  out en vdd in vss
*.iopin in
*.iopin out
*.iopin vdd
*.iopin vss
*.ipin en
XM1 vdd vg vbsh vbsh sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 vg enb vbsh vbsh sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC1 vbsh vbsl sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XM8 vbsl enb vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 vbsl vg in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 out vg in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 vs vdd vg vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 vss enb vs vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
x1 vdd en enb vss inv_lvt
.ends


* expanding   symbol:  adc/inv_lvt.sym # of pins=4
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/inv_lvt.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/inv_lvt.sch
.subckt inv_lvt  vdd in out vss
*.ipin in
*.iopin vdd
*.iopin vss
*.opin out
XM1 out in vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
