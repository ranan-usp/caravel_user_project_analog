** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/tb_switch.sch
**.subckt tb_switch
V2 net1 GND DC pulse(0 1.8 0 30p 30p 5.555n 11.11n)
V3 VIN GND DC pulse(1 1 0 12.8u 0 0.2u 13u)
V1 VDD GND 1.8
x1 net1 VOUT VIN analog_switch
C1 VOUT GND 10f m=1
**** begin user architecture code
 .lib /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice



.options acct list
.temp 25
.control
tran 10n 13u
write tb_saradc.raw
plot VIN VOUT
.endc


**** end user architecture code
**.ends

* expanding   symbol:  analog_switch.sym # of pins=3
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/analog_switch.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/analog_switch.sch
.subckt analog_switch  control OUT IN
*.ipin IN
*.ipin control
*.opin OUT
x1 net1 OUT IN control transmission_gate
x2 control net1 not
.ends


* expanding   symbol:  transmission_gate.sym # of pins=4
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/transmission_gate.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/transmission_gate.sch
.subckt transmission_gate  GP OUT IN GN
*.opin OUT
*.ipin IN
*.ipin GN
*.ipin GP
XM1 OUT GN IN GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT GP IN VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  not.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/not.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/not.sch
.subckt not  a y
*.ipin a
*.opin y
XM1 y a GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
