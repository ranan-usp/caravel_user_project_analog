** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/tb_saradc.sch
**.subckt tb_saradc Q00 Q01 Q02 Q03 Q04 Q05
*.opin Q00
*.opin Q01
*.opin Q02
*.opin Q03
*.opin Q04
*.opin Q05
x3 SW3B SW4B SW1 SW2 SW0 SW3 SW0B SW1B SW2B SW5 SW5B SW4 Q03 Q04 Q00 Q05 Q01 Q02 COMP_IN Sample CLK
+ COMP_EN my_sar_logic
V2 VIN GND DC pulse(0 1 0 12.8u 0 0.2u 13u)
V4 VDD GND 1.8
x1 Vref SW0 SW1 Sample SW3 SW0B COMP_ENB SW1B SW2 SW2B SW5B SW3B SW4 SW4B SW5 VCM VIN my_cdac
x5 CLK COMP_EN GND GND VDD VDD net2 sky130_fd_sc_hd__nor2_1
XC1 net3 GND sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
x4 COMP_EN GND GND VDD VDD COMP_ENB sky130_fd_sc_hd__inv_1
V1 CLK GND DC pulse(0 1.8 0 100p 100p 11.11n 22.22n)
V3 VCM GND 0
V5 net1 VCM 0.9
V6 net4 Vref 0.9
x2 VDD COMP_IN net3 net1 net4 net2 my_comparator
**** begin user architecture code
 .lib /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice



.options acct list
.temp 25

.tran 1n 13u
.control
save all
write tb_saradc2.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  my_sar_logic.sym # of pins=22
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_sar_logic.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_sar_logic.sch
.subckt my_sar_logic  SW3B SW4B SW1 SW2 SW0 SW3 SW0B SW1B SW2B SW5 SW5B SW4 Q03 Q04 Q00 Q05 Q01 Q02
+ COMP_IN Sample CLK COMP_EN
*.opin Sample
*.ipin COMP_IN
*.opin Q05
*.opin Q04
*.opin Q03
*.opin Q02
*.opin Q01
*.opin Q00
*.opin SW5
*.opin SW4
*.opin SW4B
*.opin SW3
*.opin SW3B
*.opin SW2
*.opin SW2B
*.opin SW1
*.opin SW1B
*.opin SW0
*.opin SW0B
*.opin SW5B
*.ipin CLK
*.opin COMP_EN
x7 SW4 GND GND VDD VDD SW4B sky130_fd_sc_hd__inv_2
x10 SW5 GND GND VDD VDD SW5B sky130_fd_sc_hd__inv_2
x13 SW3 GND GND VDD VDD SW3B sky130_fd_sc_hd__inv_2
x16 SW2 GND GND VDD VDD SW2B sky130_fd_sc_hd__inv_2
x19 SW1 GND GND VDD VDD SW1B sky130_fd_sc_hd__inv_2
x43 SW0 GND GND VDD VDD SW0B sky130_fd_sc_hd__inv_2
x47 Sample D6 5D GND GND VDD VDD SW5 sky130_fd_sc_hd__or3_1
x37 Sample D5 4D GND GND VDD VDD SW4 sky130_fd_sc_hd__or3_1
x38 Sample D4 3D GND GND VDD VDD SW3 sky130_fd_sc_hd__or3_1
x39 Sample D3 2D GND GND VDD VDD SW2 sky130_fd_sc_hd__or3_1
x40 Sample D2 1D GND GND VDD VDD SW1 sky130_fd_sc_hd__or3_1
x41 Sample D1 net1 GND GND VDD VDD SW0 sky130_fd_sc_hd__or3_1
x20 D6B 5D COMP_IN Sample my_df
x23 D5B 4D COMP_IN Sample my_df
x25 D4B 3D COMP_IN Sample my_df
x26 D3B 2D COMP_IN Sample my_df
x27 D2B 1D COMP_IN Sample my_df
x35 D1B net1 COMP_IN Sample my_df
V1 VA GND 1.8
x22 D6 GND GND VDD VDD D6B sky130_fd_sc_hd__inv_2
x24 D5 GND GND VDD VDD D5B sky130_fd_sc_hd__inv_2
x36 D4 GND GND VDD VDD D4B sky130_fd_sc_hd__inv_2
x44 D3 GND GND VDD VDD D3B sky130_fd_sc_hd__inv_2
x45 D2 GND GND VDD VDD D2B sky130_fd_sc_hd__inv_2
x46 D1 GND GND VDD VDD D1B sky130_fd_sc_hd__inv_2
x42 VA VB GND GND VDD VDD Sample sky130_fd_sc_hd__and2_0
x2 VC COMP_EN GND GND VDD VDD GND sky130_fd_sc_hd__and2_0
x4 VE VF GND GND VDD VDD D6 sky130_fd_sc_hd__and2_0
x6 VG VH GND GND VDD VDD D5 sky130_fd_sc_hd__and2_0
x9 VI VJ GND GND VDD VDD D4 sky130_fd_sc_hd__and2_0
x12 VK VL GND GND VDD VDD D3 sky130_fd_sc_hd__and2_0
x15 VM VN GND GND VDD VDD D2 sky130_fd_sc_hd__and2_0
x18 VO VP GND GND VDD VDD D1 sky130_fd_sc_hd__and2_0
x21 CLK VE VC COMP_EN mark my_df2
x28 CLK VG VE VF clear my_df2
x29 CLK VI VG VH clear my_df2
x30 CLK VK VI VJ clear my_df2
x31 CLK VM VK VL clear my_df2
x32 CLK VO VM VN clear my_df2
x33 CLK mark VO VP clear my_df2
x34 CLK GND GND VDD VDD mark2 sky130_fd_sc_hd__inv_2
x5 mark2 clear mark my_df3
x48 CLK VC VA VB clear df4
x1 clear Q05 5D my_df3
x3 clear Q04 4D my_df3
x8 clear Q03 3D my_df3
x11 clear Q02 2D my_df3
x14 clear Q01 1D my_df3
x17 clear Q00 net1 my_df3
.ends


* expanding   symbol:  my_cdac.sym # of pins=17
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_cdac.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_cdac.sch
.subckt my_cdac  Vref SW0 SW1 Sample SW3 SW0B COMP_ENB SW1B SW2 SW2B SW5B SW3B SW4 SW4B SW5 VCM VIN
*.ipin VCM
*.ipin VIN
*.ipin COMP_ENB
*.ipin Sample
*.ipin SW0
*.ipin SW0B
*.ipin SW1
*.ipin SW1B
*.ipin SW2
*.ipin SW2B
*.ipin SW3
*.ipin SW3B
*.ipin SW4
*.ipin SW4B
*.ipin SW5
*.ipin SW5B
*.opin Vref
xproblem COMP_ENB C7V VCM analog_switch
x2 Sample C7V CDACin analog_switch
x3 SW0B C6V VCM analog_switch
x4 SW0 C6V CDACin analog_switch
x5 SW1B C5V VCM analog_switch
x6 SW1 C5V CDACin analog_switch
x7 SW2B C4V VCM analog_switch
x8 SW2 C4V CDACin analog_switch
x9 SW3B C3V VCM analog_switch
x10 SW3 C3V CDACin analog_switch
x11 SW4B C2V VCM analog_switch
x12 SW4 C2V CDACin analog_switch
x13 SW5B C1V VCM analog_switch
x14 SW5 C1V CDACin analog_switch
x15 Vref C5V cap2
x16 Vref C4V cap4
x17 Vref C3V cap8
x18 Vref C2V cap16
x19 Vref C1V cap32
XC1 Vref C7V sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC2 Vref C6V sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
x1 Sample Vref GND analog_switch
x20 COMP_ENB CDACin net1 analog_switch
x21 Sample CDACin VIN analog_switch
V1 net1 GND 0
.ends


* expanding   symbol:  my_comparator.sym # of pins=6
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_comparator.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_comparator.sch
.subckt my_comparator  VDD VOUTP VOUTN VINP VINN CLK
*.ipin VDD
*.opin VOUTN
*.opin VOUTP
*.ipin CLK
*.ipin VINP
*.ipin VINN
XM2 net1 VINP net3 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=MN m=MN
XM4 net1 CLK VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=MP m=MP
**** begin user architecture code


.param MP=1
.param MN=1


**** end user architecture code
XM5 net2 CLK VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=MP m=MP
XM6 net5 net2 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=MP m=MP
XM7 net4 net1 VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=MP m=MP
XM8 VOUTP VOUTN net4 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=MP m=MP
XM9 VOUTN VOUTP net5 VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=MP m=MP
XM1 net2 VINN net3 GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=MN m=MN
XM3 net3 CLK GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=MN m=MN
XM10 net5 net2 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=MN m=MN
XM11 net4 net1 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=MN m=MN
XM12 VOUTP net1 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=MN m=MN
XM13 VOUTP VOUTN GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=MN m=MN
XM14 VOUTN net2 GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=MN m=MN
XM15 VOUTN VOUTP GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=MN m=MN
.ends


* expanding   symbol:  my_df.sym # of pins=4
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_df.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_df.sch
.subckt my_df  CLK Q D RESET
*.ipin CLK
*.ipin D
*.ipin RESET
*.opin Q
x1 RESET GND GND VDD VDD net1 sky130_fd_sc_hd__inv_1
x3 CLK D net1 GND GND VDD VDD Q sky130_fd_sc_hd__dfrtp_1
.ends


* expanding   symbol:  my_df2.sym # of pins=5
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_df2.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_df2.sch
.subckt my_df2  CLK Q D Q_N RESET
*.ipin CLK
*.ipin D
*.ipin RESET
*.opin Q
*.opin Q_N
x1 RESET GND GND VDD VDD net1 sky130_fd_sc_hd__inv_1
x2 CLK D net1 VDD GND GND VDD VDD Q Q_N sky130_fd_sc_hd__dfbbp_1
.ends


* expanding   symbol:  my_df3.sym # of pins=3
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_df3.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/my_df3.sch
.subckt my_df3  CLK Q D
*.ipin CLK
*.ipin D
*.opin Q
x1 CLK D VDD GND GND VDD VDD Q sky130_fd_sc_hd__dfrtp_1
.ends


* expanding   symbol:  df4.sym # of pins=5
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/df4.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/df4.sch
.subckt df4  CLK Q D Q_N RESET
*.ipin CLK
*.ipin D
*.ipin RESET
*.opin Q
*.opin Q_N
x2 RESET GND GND VDD VDD net1 sky130_fd_sc_hd__inv_1
x1 CLK D net1 GND GND VDD VDD Q Q_N sky130_fd_sc_hd__dfrbp_1
.ends


* expanding   symbol:  analog_switch.sym # of pins=3
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/analog_switch.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/analog_switch.sch
.subckt analog_switch  control OUT IN
*.ipin IN
*.ipin control
*.opin OUT
x1 net1 OUT IN control transmission_gate
x2 control net1 not
.ends


* expanding   symbol:  cap2.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/cap2.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/cap2.sch
.subckt cap2  out in
*.ipin in
*.opin out
XC1 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC2 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
.ends


* expanding   symbol:  cap4.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/cap4.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/cap4.sch
.subckt cap4  out in
*.ipin in
*.opin out
XC1 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC2 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC3 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC4 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
.ends


* expanding   symbol:  cap8.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/cap8.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/cap8.sch
.subckt cap8  out in
*.ipin in
*.opin out
XC1 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC2 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC3 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC4 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC5 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC6 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC7 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC8 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
.ends


* expanding   symbol:  cap16.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/cap16.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/cap16.sch
.subckt cap16  out in
*.ipin in
*.opin out
XC1 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC2 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC3 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC4 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC5 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC6 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC7 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC8 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC9 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC10 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC11 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC12 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC13 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC14 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC15 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC16 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
.ends


* expanding   symbol:  cap32.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/cap32.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/cap32.sch
.subckt cap32  out in
*.ipin in
*.opin out
XC1 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC2 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC3 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC4 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC5 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC6 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC7 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC8 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC9 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC10 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC11 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC12 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC13 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC14 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC15 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC16 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC17 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC18 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC19 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC20 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC21 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC22 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC23 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC24 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC25 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC26 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC27 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC28 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC29 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC30 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC31 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
XC32 out in sky130_fd_pr__cap_mim_m3_1 W=2 L=2.15 MF=1 m=1
.ends


* expanding   symbol:  transmission_gate.sym # of pins=4
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/transmission_gate.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/transmission_gate.sch
.subckt transmission_gate  GP OUT IN GN
*.opin OUT
*.ipin IN
*.ipin GN
*.ipin GP
XM1 OUT GN IN GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 OUT GP IN VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  not.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/not.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/not.sch
.subckt not  a y
*.ipin a
*.opin y
XM1 y a GND GND sky130_fd_pr__nfet_01v8_lvt L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 y a VDD VDD sky130_fd_pr__pfet_01v8_lvt L=0.35 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
