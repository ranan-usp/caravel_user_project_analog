** sch_path:
*+ /home/oe23ranan/caravel_user_project_analog/xschem/sub/tb/comparator/tran_comparator_trim.sch
**.subckt tran_comparator_trim
xcom vss vdd clkcc outp vp outn vn trim[4] trim[3] trim[2] trim[1] trim[0] trimb[4] trimb[3]
+ trimb[2] trimb[1] trimb[0] comparator
V1 vss GND 0
V2 vdd GND 1.4
V3 net1 GND vin
V4 vn GND vin
V10 vp net1 voff
x4 clkc vss vss vdd vdd clkcc sky130_fd_sc_hd__buf_1
xlat vdd comp net2 vss outn outp latch
Vclk1 clk GND PULSE(0 1 1e-9 1e-9 1e-9 2e-6 4e-6)
V5 cal GND 1.4
Ven en GND PULSE(0 1 0.5e-6 0.1e-6 0.1e-6 10e-6 10e-3)
V6 rstn GND 1.4
**** begin user architecture code
?

Xuut dclk drstn den dcomp dcal dvalid dres0 dres1 dres2 dres3 dres4 dres5 dres6 dres7 dsamp dctlp0
+ dctlp1 dctlp2 dctlp3 dctlp4 dctlp5 dctlp6 dctlp7 dctln0 dctln1 dctln2 dctln3 dctln4 dctln5 dctln6 dctln7
+ dtrim0 dtrim1 dtrim2 dtrim3 dtrim4 dtrimb0 dtrimb1 dtrimb2 dtrimb3 dtrimb4 dclkc sar_logic

.model adc_buff adc_bridge(in_low = 0.2 in_high=0.8)
.model dac_buff dac_bridge(out_high = 1.2)

Aad [clk rstn en comp cal] [dclk drstn den dcomp dcal] adc_buff
Ada [dctlp0 dctlp1 dctlp2 dctlp3 dctlp4 dctlp5 dctlp6 dctlp7 dctln0 dctln1 dctln2 dctln3 dctln4
+ dctln5 dctln6 dctln7 dres0 dres1 dres2 dres3 dres4 dres5 dres6 dres7 dsamp dclkc] [ctlp_0_ ctlp_1_ ctlp_2_
+ ctlp_3_ ctlp_4_ ctlp_5_ ctlp_6_ ctlp_7_ ctln_0_ ctln_1_ ctln_2_ ctln_3_ ctln_4_ ctln_5_ ctln_6_ ctln_7_
+ res0 res1 res2 res3 res4 res5 res6 res7 sample clkc] dac_buff
Ada2 [dtrim4 dtrim3 dtrim2 dtrim1 dtrim0 dtrimb4 dtrimb3 dtrimb2 dtrimb1 dtrimb0] [trim_4_ trim_3_
+ trim_2_ trim_1_ trim_0_ trimb_4_ trimb_3_ trimb_2_ trimb_1_ trimb_0_ ] dac_buff



* FET CORNERS
.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/tt.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ff.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ss.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/sf.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/fs.spice

* TT + R + C
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/tt_rmax_cmax.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/tt_rmin_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/tt_rmax_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/tt_rmin_cmax.spice

* FF + R + C
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ff_rmax_cmax.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ff_rmin_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ff_rmax_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ff_rmin_cmax.spice


* SS + R + C
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ss_rmax_cmax.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ss_rmin_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ss_rmax_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ss_rmin_cmax.spice

* SF + R + C
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/sf_rmax_cmax.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/sf_rmin_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/sf_rmax_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/sf_rmin_cmax.spice

* FS + R + C
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/fs_rmax_cmax.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/fs_rmin_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/fs_rmax_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/fs_rmin_cmax.spice

.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.ref/sky130_fd_sc_hd/spice/cells/buf/spice__buf_1.spice

**** end user architecture code
**.ends

* expanding   symbol:  sar_10b/comparator/comparator.sym # of pins=9
** sym_path:
*+ /home/oe23ranan/caravel_user_project_analog/xschem/sub/sar_10b/comparator/comparator.sym
** sch_path:
*+ /home/oe23ranan/caravel_user_project_analog/xschem/sub/sar_10b/comparator/comparator.sch
.subckt comparator  vss vdd clk outp vp outn vn trim[4] trim[3] trim[2] trim[1] trim[0] trimb[4]
+ trimb[3] trimb[2] trimb[1] trimb[0]
*.ipin vn
*.ipin vp
*.ipin clk
*.iopin vdd
*.iopin vss
*.opin outp
*.opin outn
*.ipin trim[4],trim[3],trim[2],trim[1],trim[0]
*.ipin trimb[4],trimb[3],trimb[2],trimb[1],trimb[0]
*  Mdiff -  nfet_01v8  IS MISSING !!!!
*  Minn -  nfet_01v8  IS MISSING !!!!
*  Minp -  nfet_01v8  IS MISSING !!!!
*  Ml4 -  pfet_01v8  IS MISSING !!!!
*  Ml3 -  pfet_01v8  IS MISSING !!!!
*  M3 -  pfet_01v8  IS MISSING !!!!
*  M2 -  pfet_01v8  IS MISSING !!!!
*  Ml1 -  nfet_01v8  IS MISSING !!!!
*  Ml2 -  nfet_01v8  IS MISSING !!!!
*  M4 -  pfet_01v8  IS MISSING !!!!
*  M1 -  pfet_01v8  IS MISSING !!!!
x2 in trim[4] trim[3] trim[2] trim[1] trim[0] vss trim
x3 ip trimb[4] trimb[3] trimb[2] trimb[1] trimb[0] vss trim
.ends


* expanding   symbol:  sar_10b/latch/latch.sym # of pins=6
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/sub/sar_10b/latch/latch.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/sub/sar_10b/latch/latch.sch
.subckt latch  vdd Q Qn vss R S
*.ipin S
*.ipin R
*.iopin vss
*.iopin vdd
*.opin Q
*.opin Qn
x1 vdd Qn Q vss inv_lvt
x2 vdd Q Qn vss inv_lvt
x3 vdd R net2 vss inv_lvt
x4 vdd S net1 vss inv_lvt
*  M3 -  nfet_01v8_lvt  IS MISSING !!!!
*  M1 -  nfet_01v8_lvt  IS MISSING !!!!
.ends


* expanding   symbol:  sar_10b/comparator/trim.sym # of pins=3
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/sub/sar_10b/comparator/trim.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/sub/sar_10b/comparator/trim.sch
.subckt trim  drain d[4] d[3] d[2] d[1] d[0] vss
*.iopin vss
*.ipin d[4],d[3],d[2],d[1],d[0]
*.opin drain
*  M4[7],M4[6],M4[5],M4[4],M4[3],M4[2],M4[1],M4[0] -  nfet_01v8_lvt  IS MISSING !!!!
*  M3[3],M3[2],M3[1],M3[0] -  nfet_01v8_lvt  IS MISSING !!!!
*  M2[1],M2[0] -  nfet_01v8_lvt  IS MISSING !!!!
*  M1 -  nfet_01v8_lvt  IS MISSING !!!!
*  M0 -  nfet_01v8_lvt  IS MISSING !!!!
x4[7] drain n4 trimcap
x4[6] drain n4 trimcap
x4[5] drain n4 trimcap
x4[4] drain n4 trimcap
x4[3] drain n4 trimcap
x4[2] drain n4 trimcap
x4[1] drain n4 trimcap
x4[0] drain n4 trimcap
x3[3] drain n3 trimcap
x3[2] drain n3 trimcap
x3[1] drain n3 trimcap
x3[0] drain n3 trimcap
x2[1] drain n2 trimcap
x2[0] drain n2 trimcap
x1 drain n1 trimcap
x0 drain n0 trimcap
.ends


* expanding   symbol:  logic/inv_lvt.sym # of pins=4
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/sub/logic/inv_lvt.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/sub/logic/inv_lvt.sch
.subckt inv_lvt  vdd in out vss
*.iopin vdd
*.iopin vss
*.ipin in
*.opin out
*  M1 -  nfet_01v8_lvt  IS MISSING !!!!
*  M2 -  pfet_01v8_lvt  IS MISSING !!!!
.ends


* expanding   symbol:  sar_10b/comparator/trimcap.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/sub/sar_10b/comparator/trimcap.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/sub/sar_10b/comparator/trimcap.sch
.subckt trimcap  cp cn
*.iopin cp
*.iopin cn
c0 net1 cn 2f m=1
c1 cp net1 1f m=1
.ends

.GLOBAL GND
.end
