** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/tb/cdac/tb_cdac2.sch
**.subckt tb_cdac2 aout
*.opin aout
x2 sw VGND VNB VPB VPWR swb sky130_fd_sc_hd__inv_2
V1 sw GND dummy
C1 aout net1 2.6f m=1
x1 sw VGND VNB VPB VPWR swb sky130_fd_sc_hd__inv_2
V2 sw GND d0
C2 aout net2 2.6f m=1
x3 sw VGND VNB VPB VPWR swb sky130_fd_sc_hd__inv_2
V3 sw GND d1
C3_1_ aout net3 2.6f m=1
C3_0_ aout net3 2.6f m=1
x4 sw VGND VNB VPB VPWR swb sky130_fd_sc_hd__inv_2
V4 sw GND d2
C4_3_ aout net4 2.6f m=1
C4_2_ aout net4 2.6f m=1
C4_1_ aout net4 2.6f m=1
C4_0_ aout net4 2.6f m=1
x5 sw VGND VNB VPB VPWR swb sky130_fd_sc_hd__inv_2
V5 sw GND d3
C3_7_ aout net5 2.6f m=1
C3_6_ aout net5 2.6f m=1
C3_5_ aout net5 2.6f m=1
C3_4_ aout net5 2.6f m=1
C3_3_ aout net5 2.6f m=1
C3_2_ aout net5 2.6f m=1
C3_1_ aout net5 2.6f m=1
C3_0_ aout net5 2.6f m=1
x6 sw VGND VNB VPB VPWR swb sky130_fd_sc_hd__inv_2
V6 sw GND d4
C4_15_ aout net6 2.6f m=1
C4_14_ aout net6 2.6f m=1
C4_13_ aout net6 2.6f m=1
C4_12_ aout net6 2.6f m=1
C4_11_ aout net6 2.6f m=1
C4_10_ aout net6 2.6f m=1
C4_9_ aout net6 2.6f m=1
C4_8_ aout net6 2.6f m=1
C4_7_ aout net6 2.6f m=1
C4_6_ aout net6 2.6f m=1
C4_5_ aout net6 2.6f m=1
C4_4_ aout net6 2.6f m=1
C4_3_ aout net6 2.6f m=1
C4_2_ aout net6 2.6f m=1
C4_1_ aout net6 2.6f m=1
C4_0_ aout net6 2.6f m=1
x7 sw VGND VNB VPB VPWR swb sky130_fd_sc_hd__inv_2
V7 sw GND d5
C5_31_ aout net7 2.6f m=1
C5_30_ aout net7 2.6f m=1
C5_29_ aout net7 2.6f m=1
C5_28_ aout net7 2.6f m=1
C5_27_ aout net7 2.6f m=1
C5_26_ aout net7 2.6f m=1
C5_25_ aout net7 2.6f m=1
C5_24_ aout net7 2.6f m=1
C5_23_ aout net7 2.6f m=1
C5_22_ aout net7 2.6f m=1
C5_21_ aout net7 2.6f m=1
C5_20_ aout net7 2.6f m=1
C5_19_ aout net7 2.6f m=1
C5_18_ aout net7 2.6f m=1
C5_17_ aout net7 2.6f m=1
C5_16_ aout net7 2.6f m=1
C5_15_ aout net7 2.6f m=1
C5_14_ aout net7 2.6f m=1
C5_13_ aout net7 2.6f m=1
C5_12_ aout net7 2.6f m=1
C5_11_ aout net7 2.6f m=1
C5_10_ aout net7 2.6f m=1
C5_9_ aout net7 2.6f m=1
C5_8_ aout net7 2.6f m=1
C5_7_ aout net7 2.6f m=1
C5_6_ aout net7 2.6f m=1
C5_5_ aout net7 2.6f m=1
C5_4_ aout net7 2.6f m=1
C5_3_ aout net7 2.6f m=1
C5_2_ aout net7 2.6f m=1
C5_1_ aout net7 2.6f m=1
C5_0_ aout net7 2.6f m=1
S1 net1 GND swb GND SWITCH1
S2 net1 vin sw GND SWITCH1
S3 net2 GND swb GND SWITCH1
S4 net2 vin sw GND SWITCH1
S5 net3 GND swb GND SWITCH1
S6 net3 vin sw GND SWITCH1
S7 net4 GND swb GND SWITCH1
S8 net4 vin sw GND SWITCH1
S9 net5 GND swb GND SWITCH1
S10 net5 vin sw GND SWITCH1
S11 net6 GND swb GND SWITCH1
S12 net6 vin sw GND SWITCH1
S13 net7 GND swb GND SWITCH1
S14 net7 vin sw GND SWITCH1
**** begin user architecture code
 * FET CORNERS
.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest//corners/ff.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs.spice

* TT + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmin_cmax.spice

* FF + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmin_cmax.spice


* SS + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmin_cmax.spice

* SF + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmin_cmax.spice

* FS + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmin_cmax.spice



.option wnflag=1
Vin vin 0 PULSE 0 1 0 12.8u 0 0.2u 13u

.control
save all
tran 13u 1u

.param dummy=1
.param d5=0
.param d4=1
.param d3=1
.param d2=1
.param d1=1
.param d0=1



op
write test_cdac.raw
.endc




.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_2.spice
**** end user architecture code
**.ends
.GLOBAL GND
.end
