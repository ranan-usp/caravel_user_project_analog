** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/tb/cdac/tb_cdac3.sch
**.subckt tb_cdac3
V1 sw GND dummy
V2 sw1 GND d0
V3 sw2 GND d1
V4 sw3 GND d2
V5 sw4 GND d3
V6 sw5 GND d4
V7 sw6 GND d5
x10 in_dummy swbd vdd GND vss my_passgate
x11 in_dummy sw vdd vin vss my_passgate
x12 in1 swb1 vdd GND vss my_passgate
x13 in1 sw1 vdd vin vss my_passgate
x14 in2 swb2 vdd GND vss my_passgate
x15 in2 sw2 vdd vin vss my_passgate
x16 in3 swb3 vdd GND vss my_passgate
x17 in3 sw3 vdd vin vss my_passgate
x18 in4 swb4 vdd GND vss my_passgate
x19 in4 sw4 vdd vin vss my_passgate
x20 in5 swb5 vdd GND vss my_passgate
x21 in5 sw5 vdd vin vss my_passgate
x22 in6 swb6 vdd GND vss my_passgate
x23 in6 sw6 vdd vin vss my_passgate
x7 sw6 vss vss vdd vdd swb6 sky130_fd_sc_hd__inv_2
x1 sw5 vss vss vdd vdd swb5 sky130_fd_sc_hd__inv_2
x2 sw4 vss vss vdd vdd swb4 sky130_fd_sc_hd__inv_2
x3 sw3 vss vss vdd vdd swb3 sky130_fd_sc_hd__inv_2
x4 sw2 vss vss vdd vdd swb2 sky130_fd_sc_hd__inv_2
x5 sw1 vss vss vdd vdd swb1 sky130_fd_sc_hd__inv_2
x6 sw vss vss vdd vdd swbd sky130_fd_sc_hd__inv_2
R7 dd0 ddummy para m=1
R1 dd1 dd0 para m=1
R2 dd2 dd1 para m=1
R3 dd3 dd2 para m=1
R4 dd4 dd3 para m=1
R5 output dd4 para m=1
R_para_dummy in_dummy in_dummy_dash 5 m=1
R_para1 in1 in1_dash 5 m=1
R_para2 in2 in2_dash 5 m=1
R_para3 in3 in3_dash 5 m=1
R_para4 in4 in4_dash 5 m=1
R_para5 in5 in5_dash 5 m=1
R_para6 in6 in6_dash 5 m=1
CP0 ddummy in_dummy_dash 1p m=1
CP1 dd0 in1_dash 1p m=1
CP2 dd1 in2_dash 1p m=1
CP3 dd2 in3_dash 1p m=1
CP4 dd3 in4_dash 1p m=1
CP5 dd4 in5_dash 1p m=1
CP6 output in6_dash 1p m=1
**** begin user architecture code
 * FET CORNERS
.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs.spice

* TT + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmin_cmax.spice

* FF + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmin_cmax.spice


* SS + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmin_cmax.spice

* SF + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmin_cmax.spice

* FS + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmin_cmax.spice



.option wnflag=1
.option plotwinsize=0
Vin vin 0 dc PULSE(0 1 0 12.8u 0 0.2u 13u)
*Vin vin 0 1.8
VDD vdd 0 1.8
VSS vss 0 0

.param dummy=0
.param d5=1
.param d4=0
.param d3=0
.param d2=0
.param d1=0
.param d0=0
.param para=5

.control
save all
tran 1u 13u

meas tran output find v(d5) at=13u

wrdata out output
print output
.endc




.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_2.spice
**** end user architecture code
**.ends

* expanding   symbol:  switches/my_passgate.sym # of pins=5
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/switches/my_passgate.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/switches/my_passgate.sch
.subckt my_passgate  out en vdd in vss
*.iopin out
*.ipin en
*.iopin vss
*.iopin vdd
*.iopin in
x2 vdd en enb vss inv_lvt
x1 vdd enb en_buf vss inv_lvt
XMSN out en_buf in vss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMSP in enb out vdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  logic/inv_lvt.sym # of pins=4
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/logic/inv_lvt.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/logic/inv_lvt.sch
.subckt inv_lvt  vdd in out vss
*.iopin vdd
*.iopin vss
*.ipin in
*.opin out
XM1 out in vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
