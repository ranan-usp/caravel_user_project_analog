** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/sarlogic.sch
**.subckt sarlogic comp cal en clk valid rstn
*+ result[9],result[8],result[7],result[6],result[5],result[4],result[3],result[2],result[1],result[0] trimb[4],trimb[3],trimb[2],trimb[1],trimb[0] trim[4],trim[3],trim[2],trim[1],trim[0] clkc sample
*+ ctlp[9],ctlp[8],ctlp[7],ctlp[6],ctlp[5],ctlp[4],ctlp[3],ctlp[2],ctlp[1],ctlp[0] ctln[9],ctln[8],ctln[7],ctln[6],ctln[5],ctln[4],ctln[3],ctln[2],ctln[1],ctln[0] dvdd dvss
*.ipin comp
*.ipin cal
*.ipin en
*.ipin clk
*.ipin valid
*.ipin rstn
*.ipin
*+ result[9],result[8],result[7],result[6],result[5],result[4],result[3],result[2],result[1],result[0]
*.opin trimb[4],trimb[3],trimb[2],trimb[1],trimb[0]
*.opin trim[4],trim[3],trim[2],trim[1],trim[0]
*.opin clkc
*.opin sample
*.opin ctlp[9],ctlp[8],ctlp[7],ctlp[6],ctlp[5],ctlp[4],ctlp[3],ctlp[2],ctlp[1],ctlp[0]
*.opin ctln[9],ctln[8],ctln[7],ctln[6],ctln[5],ctln[4],ctln[3],ctln[2],ctln[1],ctln[0]
*.iopin dvdd
*.iopin dvss
**** begin user architecture code
.include /home/oe23ranan/caravel_user_project_analog/xschem/adc/cmos_cells_digital.sp
.include /home/oe23ranan/caravel_user_project_analog/xschem/adc/sarlogic.sp

**** end user architecture code
**.ends
.end
