** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/6bit_saradc.sch
**.subckt 6bit_saradc vdd vss dvdd dvss vinp vinn clk Q[5],Q[4],Q[3],Q[2],Q[1],Q[0]
*.iopin vdd
*.iopin vss
*.iopin dvdd
*.iopin dvss
*.ipin vinp
*.ipin vinn
*.ipin clk
*.opin Q[5],Q[4],Q[3],Q[2],Q[1],Q[0]
x3 vss vdd clkc net3 net1 net4 net2 comp
x4 vdd net6 net5 vss net4 net3 latch
x5 dvdd dvss clk net6 sample clkc Q[5] Q[4] Q[3] Q[2] Q[1] Q[0] ctrl[5] ctrl[4] ctrl[3] ctrl[2]
+ ctrl[1] ctrl[0] ctrlb[5] ctrlb[4] ctrlb[3] ctrlb[2] ctrlb[1] ctrlb[0] my_sar_logic
x1 net1 sample vdd vss vinp ctrl[5] ctrl[4] ctrl[3] ctrl[2] ctrl[1] ctrl[0] vdd dac
x2 net2 sample vdd vss vinn ctrlb[5] ctrlb[4] ctrlb[3] ctrlb[2] ctrlb[1] ctrlb[0] vss dac
**.ends

* expanding   symbol:  adc/comp.sym # of pins=7
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/comp.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/comp.sch
.subckt comp  vss vdd clk outp vp outn vn
*.ipin vn
*.ipin vp
*.ipin clk
*.iopin vdd
*.iopin vss
*.opin outp
*.opin outn
XMl1 outn outp net1 vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMl2 outp outn net2 vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMinp net2 vp diff vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMinn net1 vn diff vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMdiff diff clk vss vss sky130_fd_pr__nfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 outn clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 outp outn vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 outn outp vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 outp clk vdd vdd sky130_fd_pr__pfet_01v8 L=0.3 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc/latch.sym # of pins=6
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/latch.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/latch.sch
.subckt latch  vdd Q Qn vss R S
*.ipin S
*.ipin R
*.iopin vss
*.iopin vdd
*.opin Q
*.opin Qn
x1 vdd Qn Q vss inv_lvt
x2 vdd Q Qn vss inv_lvt
x3 vdd R net2 vss inv_lvt
x4 vdd S net1 vss inv_lvt
XM1 Qn net1 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Q net2 vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc/my_sar_logic.sym # of pins=9
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/my_sar_logic.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/my_sar_logic.sch
.subckt my_sar_logic  dvdd dvss CLK COMP_IN Sample clkc Q[5] Q[4] Q[3] Q[2] Q[1] Q[0] SW[5] SW[4]
+ SW[3] SW[2] SW[1] SW[0] SWB[5] SWB[4] SWB[3] SWB[2] SWB[1] SWB[0]
*.opin Sample
*.ipin COMP_IN
*.ipin CLK
*.opin clkc
*.opin Q[5],Q[4],Q[3],Q[2],Q[1],Q[0]
*.opin SW[5],SW[4],SW[3],SW[2],SW[1],SW[0]
*.opin SWB[5],SWB[4],SWB[3],SWB[2],SWB[1],SWB[0]
*.iopin dvss
*.iopin dvdd
x41 Sample D1 net2 avss dvss dvdd dvdd SW[0] sky130_fd_sc_hd__or3_1
x46 D1 dvss dvss dvdd dvdd D1B sky130_fd_sc_hd__inv_2
x22 D2 dvss dvss dvdd dvdd D2B sky130_fd_sc_hd__inv_2
x24 D3 dvss dvss dvdd dvdd D3B sky130_fd_sc_hd__inv_2
x34 D4 dvss dvss dvdd dvdd D4B sky130_fd_sc_hd__inv_2
x36 D5 dvss dvss dvdd dvdd D5B sky130_fd_sc_hd__inv_2
x44 D6 dvss dvss dvdd dvdd D6B sky130_fd_sc_hd__inv_2
x45 CLK dvss dvss dvdd dvdd mark2 sky130_fd_sc_hd__inv_2
x49 CLK COMP_EN dvss dvss dvdd Vdvdd clkc sky130_fd_sc_hd__nor2_1
x1 CLK VC dvdd VB net1 mydf
x3 CLK VE VC COMP_EN mark mydf
x5 CLK VG VE VF net1 mydf
x8 CLK VI VG VH net1 mydf
x11 CLK VK VI VJ net1 mydf
x14 CLK VM VK VL net1 mydf
x17 CLK VO VM VN net1 mydf
x20 CLK mark VO VP net1 mydf
x23 D6B 5D COMP_IN net5 Sample mydf
x25 D5B 4D COMP_IN net6 Sample mydf
x26 D4B 3D COMP_IN net7 Sample mydf
x27 D3B 2D COMP_IN net8 Sample mydf
x28 D2B 1D COMP_IN net9 Sample mydf
x29 D1B net2 COMP_IN net10 Sample mydf
x30 mark2 net1 mark net11 net4 mydf
x31 net1 Q[5] 5D net12 net13 mydf
x32 net1 Q[4] 4D net14 net15 mydf
x33 net1 Q[3] 3D net16 net17 mydf
x35 net1 Q[2] 2D net18 net19 mydf
x48 net1 Q[1] 1D net20 net21 mydf
x50 net1 Q[0] net2 net22 net23 mydf
x18 VM VN dvss dvss dvdd dvdd D2 sky130_fd_sc_hd__and2_0
x2 VO VP dvss dvss dvdd dvdd D1 sky130_fd_sc_hd__and2_0
x4 VI VJ dvss dvss dvdd dvdd D4 sky130_fd_sc_hd__and2_0
x6 VK VL dvss dvss dvdd dvdd D3 sky130_fd_sc_hd__and2_0
x9 VE VF dvss dvss dvdd dvdd D6 sky130_fd_sc_hd__and2_0
x12 VG VH dvss dvss dvdd dvdd D5 sky130_fd_sc_hd__and2_0
x15 dvdd VB dvss dvss dvdd dvdd Sample sky130_fd_sc_hd__and2_0
x42 VC COMP_EN dvss dvss dvdd dvdd net3 sky130_fd_sc_hd__and2_0
x7 SW[0] dvss dvss dvdd dvdd SWB[0] sky130_fd_sc_hd__inv_2
x10 SW[1] dvss dvss dvdd dvdd SWB[1] sky130_fd_sc_hd__inv_2
x13 SW[2] dvss dvss dvdd dvdd SWB[2] sky130_fd_sc_hd__inv_2
x16 SW[3] dvss dvss dvdd dvdd SWB[3] sky130_fd_sc_hd__inv_2
x19 SW[4] dvss dvss dvdd dvdd SWB[4] sky130_fd_sc_hd__inv_2
x43 SW[5] dvss dvss dvdd dvdd SWB[5] sky130_fd_sc_hd__inv_2
x37 Sample D2 1D avss dvss dvdd dvdd SW[1] sky130_fd_sc_hd__or3_1
x38 Sample D3 2D avss dvss dvdd dvdd SW[2] sky130_fd_sc_hd__or3_1
x39 Sample D4 3D avss dvss dvdd dvdd SW[3] sky130_fd_sc_hd__or3_1
x40 Sample D5 4D avss dvss dvdd dvdd SW[4] sky130_fd_sc_hd__or3_1
x47 Sample D6 5D avss dvss dvdd dvdd SW[5] sky130_fd_sc_hd__or3_1
.ends


* expanding   symbol:  adc/dac.sym # of pins=7
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/dac.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/dac.sch
.subckt dac  out sample vdd vss vin ctrl[5] ctrl[4] ctrl[3] ctrl[2] ctrl[1] ctrl[0] dum
*.opin out
*.ipin vin
*.ipin sample
*.ipin ctrl[5],ctrl[4],ctrl[3],ctrl[2],ctrl[1],ctrl[0]
*.ipin dum
*.iopin vdd
*.iopin vss
x1 out ctrl[0] net5 net4 net2 dum net3 net1 carry
x2 out sample vdd vin vss bootstrapped_sw_hv
xi4 ctrl[5] vss vss vdd vdd net5 sky130_fd_sc_hd__inv_2
xi5 ctrl[4] vss vss vdd vdd net4 sky130_fd_sc_hd__inv_2
xi6 ctrl[3] vss vss vdd vdd net3 sky130_fd_sc_hd__inv_2
xi7 ctrl[2] vss vss vdd vdd net2 sky130_fd_sc_hd__inv_2
xi9 ctrl[1] vss vss vdd vdd net1 sky130_fd_sc_hd__inv_2
.ends


* expanding   symbol:  adc/inv_lvt.sym # of pins=4
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/inv_lvt.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/inv_lvt.sch
.subckt inv_lvt  vdd in out vss
*.ipin in
*.iopin vdd
*.iopin vss
*.opin out
XM1 out in vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  adc/mydf.sym # of pins=5
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/mydf.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/mydf.sch
.subckt mydf  CLK Q D Q_N RESET
*.ipin CLK
*.ipin D
*.ipin RESET
*.opin Q
*.opin Q_N
x50 CLK D net1 dvss dvss dvdd dvdd Q Q_N sky130_fd_sc_hd__dfrbp_1
x1 RESET dvss dvss dvdd dvdd net1 sky130_fd_sc_hd__inv_1
.ends


* expanding   symbol:  adc/carry.sym # of pins=8
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/carry.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/carry.sch
.subckt carry  top n0 n5 n4 n2 ndum n3 n1
*.iopin n5
*.iopin n4
*.iopin n3
*.iopin n2
*.iopin n1
*.iopin n0
*.iopin ndum
*.iopin top
xc0 top n0 unit_cap
xcdum top ndum unit_cap
xc1[1] top n1 unit_cap
xc1[0] top n1 unit_cap
xc2[3] top n2 unit_cap
xc2[2] top n2 unit_cap
xc2[1] top n2 unit_cap
xc2[0] top n2 unit_cap
xc3[7] top n3 unit_cap
xc3[6] top n3 unit_cap
xc3[5] top n3 unit_cap
xc3[4] top n3 unit_cap
xc3[3] top n3 unit_cap
xc3[2] top n3 unit_cap
xc3[1] top n3 unit_cap
xc3[0] top n3 unit_cap
xc4[15] top n4 unit_cap
xc4[14] top n4 unit_cap
xc4[13] top n4 unit_cap
xc4[12] top n4 unit_cap
xc4[11] top n4 unit_cap
xc4[10] top n4 unit_cap
xc4[9] top n4 unit_cap
xc4[8] top n4 unit_cap
xc4[7] top n4 unit_cap
xc4[6] top n4 unit_cap
xc4[5] top n4 unit_cap
xc4[4] top n4 unit_cap
xc4[3] top n4 unit_cap
xc4[2] top n4 unit_cap
xc4[1] top n4 unit_cap
xc4[0] top n4 unit_cap
xc5[31] top n5 unit_cap
xc5[30] top n5 unit_cap
xc5[29] top n5 unit_cap
xc5[28] top n5 unit_cap
xc5[27] top n5 unit_cap
xc5[26] top n5 unit_cap
xc5[25] top n5 unit_cap
xc5[24] top n5 unit_cap
xc5[23] top n5 unit_cap
xc5[22] top n5 unit_cap
xc5[21] top n5 unit_cap
xc5[20] top n5 unit_cap
xc5[19] top n5 unit_cap
xc5[18] top n5 unit_cap
xc5[17] top n5 unit_cap
xc5[16] top n5 unit_cap
xc5[15] top n5 unit_cap
xc5[14] top n5 unit_cap
xc5[13] top n5 unit_cap
xc5[12] top n5 unit_cap
xc5[11] top n5 unit_cap
xc5[10] top n5 unit_cap
xc5[9] top n5 unit_cap
xc5[8] top n5 unit_cap
xc5[7] top n5 unit_cap
xc5[6] top n5 unit_cap
xc5[5] top n5 unit_cap
xc5[4] top n5 unit_cap
xc5[3] top n5 unit_cap
xc5[2] top n5 unit_cap
xc5[1] top n5 unit_cap
xc5[0] top n5 unit_cap
.ends


* expanding   symbol:  adc/bootstrapped_sw_hv.sym # of pins=5
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/bootstrapped_sw_hv.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/bootstrapped_sw_hv.sch
.subckt bootstrapped_sw_hv  out en vdd in vss
*.iopin in
*.iopin out
*.iopin vdd
*.iopin vss
*.ipin en
XM1 vdd vg vbsh vbsh sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 vg enb vbsh vbsh sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XC1 vbsh vbsl sky130_fd_pr__cap_mim_m3_1 W=5 L=5 MF=1 m=1
XM8 vbsl enb vss vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 vbsl vg in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 out vg in vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 vs vdd vg vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 vss enb vs vss sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
x1 vdd en enb vss inv_lvt
.ends


* expanding   symbol:  adc/unit_cap.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/unit_cap.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/unit_cap.sch
.subckt unit_cap  cp cn
*.iopin cp
*.iopin cn
C1 cp cn 2.6f m=1
.ends

.end
