** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/tb/cdac/tb_cdac2.sch
**.subckt tb_cdac2
V1 sw GND dummy
V2 sw1 GND d0
V3 sw2 GND d1
V4 sw3 GND d2
V5 sw4 GND d3
V6 sw5 GND d4
V7 sw6 GND d5
x9 d0 in0 unitcap
x10_1_ d1 in1 unitcap
x10_0_ d1 in1 unitcap
x11_3_ d2 in2 unitcap
x11_2_ d2 in2 unitcap
x11_1_ d2 in2 unitcap
x11_0_ d2 in2 unitcap
x12_7_ d3 in3 unitcap
x12_6_ d3 in3 unitcap
x12_5_ d3 in3 unitcap
x12_4_ d3 in3 unitcap
x12_3_ d3 in3 unitcap
x12_2_ d3 in3 unitcap
x12_1_ d3 in3 unitcap
x12_0_ d3 in3 unitcap
x13_15_ d4 in4 unitcap
x13_14_ d4 in4 unitcap
x13_13_ d4 in4 unitcap
x13_12_ d4 in4 unitcap
x13_11_ d4 in4 unitcap
x13_10_ d4 in4 unitcap
x13_9_ d4 in4 unitcap
x13_8_ d4 in4 unitcap
x13_7_ d4 in4 unitcap
x13_6_ d4 in4 unitcap
x13_5_ d4 in4 unitcap
x13_4_ d4 in4 unitcap
x13_3_ d4 in4 unitcap
x13_2_ d4 in4 unitcap
x13_1_ d4 in4 unitcap
x13_0_ d4 in4 unitcap
x14_31_ d5 in5 unitcap
x14_30_ d5 in5 unitcap
x14_29_ d5 in5 unitcap
x14_28_ d5 in5 unitcap
x14_27_ d5 in5 unitcap
x14_26_ d5 in5 unitcap
x14_25_ d5 in5 unitcap
x14_24_ d5 in5 unitcap
x14_23_ d5 in5 unitcap
x14_22_ d5 in5 unitcap
x14_21_ d5 in5 unitcap
x14_20_ d5 in5 unitcap
x14_19_ d5 in5 unitcap
x14_18_ d5 in5 unitcap
x14_17_ d5 in5 unitcap
x14_16_ d5 in5 unitcap
x14_15_ d5 in5 unitcap
x14_14_ d5 in5 unitcap
x14_13_ d5 in5 unitcap
x14_12_ d5 in5 unitcap
x14_11_ d5 in5 unitcap
x14_10_ d5 in5 unitcap
x14_9_ d5 in5 unitcap
x14_8_ d5 in5 unitcap
x14_7_ d5 in5 unitcap
x14_6_ d5 in5 unitcap
x14_5_ d5 in5 unitcap
x14_4_ d5 in5 unitcap
x14_3_ d5 in5 unitcap
x14_2_ d5 in5 unitcap
x14_1_ d5 in5 unitcap
x14_0_ d5 in5 unitcap
x10 in_dummy swbd vdd GND vss my_passgate
x11 in_dummy sw vdd vin vss my_passgate
x12 in0 swb1 vdd GND vss my_passgate
x13 in0 sw1 vdd vin vss my_passgate
x14 in1 swb2 vdd GND vss my_passgate
x15 in1 sw2 vdd vin vss my_passgate
x16 in2 swb3 vdd GND vss my_passgate
x17 in2 sw3 vdd vin vss my_passgate
x18 in3 swb4 vdd GND vss my_passgate
x19 in3 sw4 vdd vin vss my_passgate
x20 in4 swb5 vdd GND vss my_passgate
x21 in4 sw5 vdd vin vss my_passgate
x22 in5 swb6 vdd GND vss my_passgate
x23 in5 sw6 vdd vin vss my_passgate
x7 sw6 vss vss vdd vdd swb6 sky130_fd_sc_hd__inv_2
x1 sw5 vss vss vdd vdd swb5 sky130_fd_sc_hd__inv_2
x2 sw4 vss vss vdd vdd swb4 sky130_fd_sc_hd__inv_2
x3 sw3 vss vss vdd vdd swb3 sky130_fd_sc_hd__inv_2
x4 sw2 vss vss vdd vdd swb2 sky130_fd_sc_hd__inv_2
x5 sw1 vss vss vdd vdd swb1 sky130_fd_sc_hd__inv_2
x6 sw vss vss vdd vdd swbd sky130_fd_sc_hd__inv_2
x8 dummy in_dummy unitcap
R7 d0 dummy para m=1
R1 d1 d0 para m=1
R2 d2 d1 para m=1
R3 d3 d2 para m=1
R4 d4 d3 para m=1
R5 d5 d4 para m=1
**** begin user architecture code
 * FET CORNERS
.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/models/corners/tt.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs.spice

* TT + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/tt_rmin_cmax.spice

* FF + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ff_rmin_cmax.spice


* SS + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/ss_rmin_cmax.spice

* SF + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/sf_rmin_cmax.spice

* FS + R + C
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmax_cmax.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmin_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmax_cmin.spice
*.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_pr_ngspice/latest/corners/fs_rmin_cmax.spice



.option wnflag=1
.option plotwinsize=0
Vin vin 0 dc PULSE(0 1 0 12.8u 0 0.2u 13u)
*Vin vin 0 1.8
VDD vdd 0 1.8
VSS vss 0 0

.param dummy=0
.param d5=1
.param d4=0
.param d3=0
.param d2=0
.param d1=0
.param d0=0
.param para=5

.control
save all
tran 1u 13u

meas tran output find v(d5) at=13u

wrdata out output
print output
.endc




.include /home/oe23ranan/skywater/skywater-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_2.spice
**** end user architecture code
**.ends

* expanding   symbol:  sar_10b/unitcap/unitcap.sym # of pins=2
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/sar_10b/unitcap/unitcap.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/sar_10b/unitcap/unitcap.sch
.subckt unitcap  cp cn
*.iopin cp
*.iopin cn
C1 cp cn 2.6f m=1
.ends


* expanding   symbol:  switches/my_passgate.sym # of pins=5
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/switches/my_passgate.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/switches/my_passgate.sch
.subckt my_passgate  out en vdd in vss
*.iopin out
*.ipin en
*.iopin vss
*.iopin vdd
*.iopin in
x2 vdd en enb vss inv_lvt
x1 vdd enb en_buf vss inv_lvt
XMSN out en_buf in vss sky130_fd_pr__nfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XMSP in enb out vdd sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  logic/inv_lvt.sym # of pins=4
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/logic/inv_lvt.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/logic/inv_lvt.sch
.subckt inv_lvt  vdd in out vss
*.iopin vdd
*.iopin vss
*.ipin in
*.opin out
XM1 out in vss vss sky130_fd_pr__nfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out in vdd vdd sky130_fd_pr__pfet_01v8_lvt L=0.4 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
