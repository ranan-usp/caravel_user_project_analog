** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/tb_sarlogic.sch
**.subckt tb_sarlogic
x1 vdd vss trimb[4] trimb[3] trimb[2] trimb[1] trimb[0] comp cal trim[4] trim[3] trim[2] trim[1]
+ trim[0] en clk clkc sample result[9] result[8] result[7] result[6] result[5] result[4] result[3] result[2]
+ result[1] result[0] ctlp[9] ctlp[8] ctlp[7] ctlp[6] ctlp[5] ctlp[4] ctlp[3] ctlp[2] ctlp[1] ctlp[0] valid
+ ctln[9] ctln[8] ctln[7] ctln[6] ctln[5] ctln[4] ctln[3] ctln[2] ctln[1] ctln[0] rstn sarlogic
Vcomp comp GND DC 0 PULSE(0 {vdd} 40e-6 1e-9 1e-9 99e-6 100e-6)
Vrstn rstn GND DC 0 PULSE(0 1.2 10e-6 1e-9 1e-9 99e-6 100e-6)
Vclk clk GND DC 0 PULSE(0 1.2 10e-6 1e-9 1e-9 99e-6 100e-6)
V3 cal GND 0
V4 en GND {vdd}
V1 vdd GND {vdd}
V2 vss GND 0
**** begin user architecture code
 *.options method = trap
*.options gmin   = 1e-12
*.options abstol = 1e-8
*.options chtol  = 1e-18
*.options reltol = 0.01
*.options vntol  = 0.1e-6

*.options rshunt = 10e-12

.param MC_SWITCH=0

.ic v(valid)=0
.ic v(sample)=0
.ic v(clkc)=0

.ic v(trim_0_)=0
.ic v(trim_1_)=0
.ic v(trim_2_)=0
.ic v(trim_3_)=0
.ic v(trim_4_)=0
.ic v(trimb_0_)=0
.ic v(trimb_1_)=0
.ic v(trimb_2_)=0
.ic v(trimb_3_)=0
.ic v(trimb_4_)=0


.ic v(result_0_)=0
.ic v(result_1_)=0
.ic v(result_2_)=0
.ic v(result_3_)=0
.ic v(result_4_)=0
.ic v(result_5_)=0
.ic v(result_6_)=0
.ic v(result_7_)=0
.ic v(result_8_)=0
.ic v(result_9_)=0

.ic v(ctlp_0_)=0
.ic v(ctlp_1_)=0
.ic v(ctlp_2_)=0
.ic v(ctlp_3_)=0
.ic v(ctlp_4_)=0
.ic v(ctlp_5_)=0
.ic v(ctlp_6_)=0
.ic v(ctlp_7_)=0
.ic v(ctlp_8_)=0
.ic v(ctlp_9_)=0

.ic v(ctln_0_)=0
.ic v(ctln_1_)=0
.ic v(ctln_2_)=0
.ic v(ctln_3_)=0
.ic v(ctln_4_)=0
.ic v(ctln_5_)=0
.ic v(ctln_6_)=0
.ic v(ctln_7_)=0
.ic v(ctln_8_)=0
.ic v(ctln_9_)=0

.include /home/oe23ranan/caravel_user_project_analog/xschem/adc/sarlogic.ext.spice

.param vdd=1.2

*.tran 100e-9 68e-6
.tran 100e-9 68e-6 uic

.control
run

echo Simulation Finished
echo -------------------
shell date
echo -------------------

.endc

 * FET CORNERS
.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/tt.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ff.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ss.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/sf.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/fs.spice

* TT + R + C
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/tt_rmax_cmax.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/tt_rmin_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/tt_rmax_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/tt_rmin_cmax.spice

* FF + R + C
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ff_rmax_cmax.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ff_rmin_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ff_rmax_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ff_rmin_cmax.spice


* SS + R + C
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ss_rmax_cmax.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ss_rmin_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ss_rmax_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/ss_rmin_cmax.spice

* SF + R + C
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/sf_rmax_cmax.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/sf_rmin_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/sf_rmax_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/sf_rmin_cmax.spice

* FS + R + C
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/fs_rmax_cmax.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/fs_rmin_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/fs_rmax_cmin.spice
*.include /home/oe23ranan/pdk/volare/sky130/versions/41c0908b47130d5675ff8484255b43f66463a7d6/sky130A/libs.tech/ngspice/corners/fs_rmin_cmax.spice

.include /pdk/open_pdks/sources/sky130-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_4.spice
.include /pdk/open_pdks/sources/sky130-pdk/libraries/sky130_fd_sc_hd/latest/cells/decap/sky130_fd_sc_hd__decap_8.spice
.include /pdk/open_pdks/sources/sky130-pdk/libraries/sky130_fd_sc_hd/latest/cells/decap/sky130_fd_sc_hd__decap_3.spice
.include /pdk/open_pdks/sources/sky130-pdk/libraries/sky130_fd_sc_hd/latest/cells/buf/sky130_fd_sc_hd__buf_1.spice
.include /pdk/open_pdks/sources/sky130-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_1.spice
.include /pdk/open_pdks/sources/sky130-pdk/libraries/sky130_fd_sc_hd/latest/cells/inv/sky130_fd_sc_hd__inv_2.spice
.include /pdk/open_pdks/sources/sky130-pdk/libraries/sky130_fd_sc_hd/latest/cells/tap/sky130_fd_sc_hd__tap_2.spice
**** end user architecture code
**.ends

* expanding   symbol:  adc/sarlogic.sym # of pins=15
** sym_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/sarlogic.sym
** sch_path: /home/oe23ranan/caravel_user_project_analog/xschem/adc/sarlogic.sch
.subckt sarlogic  dvdd dvss trimb[4] trimb[3] trimb[2] trimb[1] trimb[0] comp cal trim[4] trim[3]
+ trim[2] trim[1] trim[0] en clk clkc sample result[9] result[8] result[7] result[6] result[5] result[4]
+ result[3] result[2] result[1] result[0] ctlp[9] ctlp[8] ctlp[7] ctlp[6] ctlp[5] ctlp[4] ctlp[3] ctlp[2]
+ ctlp[1] ctlp[0] valid ctln[9] ctln[8] ctln[7] ctln[6] ctln[5] ctln[4] ctln[3] ctln[2] ctln[1] ctln[0] rstn
*.ipin comp
*.ipin cal
*.ipin en
*.ipin clk
*.ipin valid
*.ipin rstn
*.ipin
*+ result[9],result[8],result[7],result[6],result[5],result[4],result[3],result[2],result[1],result[0]
*.opin trimb[4],trimb[3],trimb[2],trimb[1],trimb[0]
*.opin trim[4],trim[3],trim[2],trim[1],trim[0]
*.opin clkc
*.opin sample
*.opin ctlp[9],ctlp[8],ctlp[7],ctlp[6],ctlp[5],ctlp[4],ctlp[3],ctlp[2],ctlp[1],ctlp[0]
*.opin ctln[9],ctln[8],ctln[7],ctln[6],ctln[5],ctln[4],ctln[3],ctln[2],ctln[1],ctln[0]
*.iopin dvdd
*.iopin dvss
**** begin user architecture code
.include /home/oe23ranan/caravel_user_project_analog/xschem/adc/cmos_cells_digital.sp
.include /home/oe23ranan/caravel_user_project_analog/xschem/adc/sarlogic.sp

**** end user architecture code
.ends

.GLOBAL GND
.end
